magic
tech scmos
timestamp 1669647866
<< metal1 >>
rect -686 1352 3999 1367
rect -686 198 -671 1352
rect -54 987 272 990
rect -54 985 629 987
rect 914 985 918 987
rect -54 983 918 985
rect -54 890 -50 983
rect 268 887 272 983
rect -72 686 -68 795
rect 44 736 48 863
rect 0 732 48 736
rect 79 742 93 744
rect 366 742 370 862
rect 79 738 370 742
rect 0 714 7 732
rect 79 717 93 738
rect 79 716 88 717
rect -467 682 -68 686
rect -2857 196 -520 198
rect -467 196 -463 682
rect 412 543 416 983
rect 625 981 918 983
rect 625 887 629 981
rect 914 887 918 981
rect 3283 956 3820 961
rect 1627 947 2034 950
rect 1627 945 2368 947
rect 730 857 740 861
rect 730 660 734 857
rect 1008 724 1012 863
rect 793 720 1012 724
rect 793 670 797 720
rect 717 656 734 660
rect 1627 549 1632 945
rect 2029 942 2368 945
rect 2029 886 2034 942
rect 2363 887 2368 942
rect 2153 760 2157 860
rect 2153 756 2179 760
rect 2175 725 2179 756
rect 2461 754 2465 861
rect 2276 750 2465 754
rect 2276 721 2280 750
rect 3283 552 3288 956
rect 3522 911 3527 956
rect 3815 913 3820 956
rect 3625 800 3629 881
rect 3680 822 3710 837
rect 3680 809 3695 822
rect 3625 796 3642 800
rect 3638 744 3642 796
rect 3680 794 3708 809
rect 3693 778 3708 794
rect 3693 763 3726 778
rect 3711 753 3726 763
rect 3984 753 3999 1352
rect 3711 738 3999 753
rect 4187 888 5704 925
rect 4187 549 4224 888
rect -2857 192 -457 196
rect -2857 191 -520 192
rect -2855 -2665 -2850 191
rect -467 -71 -463 192
rect 451 -71 455 208
rect -467 -75 455 -71
rect 1750 -182 1782 139
rect -805 -214 1782 -182
rect -805 -1421 -773 -214
rect 3337 -399 3384 163
rect -844 -1453 -773 -1421
rect 302 -446 3384 -399
rect -844 -2004 -812 -1453
rect -374 -1752 -370 -1591
rect -746 -1756 -370 -1752
rect -746 -1762 -741 -1756
rect -745 -1977 -741 -1762
rect 52 -1973 56 -1884
rect -99 -1977 56 -1973
rect -745 -1980 -733 -1977
rect -745 -1981 -730 -1980
rect -741 -1984 -730 -1981
rect -99 -2038 -95 -1977
rect 302 -2002 349 -446
rect 4808 -602 4842 185
rect 1544 -636 4842 -602
rect 923 -1698 1351 -1694
rect 1347 -1952 1351 -1698
rect 1544 -1950 1578 -636
rect 5098 -1578 5129 185
rect 2120 -1610 2150 -1606
rect 2146 -1658 2150 -1610
rect 2863 -1609 5129 -1578
rect 2146 -1662 2693 -1658
rect 1346 -1962 1369 -1952
rect 1347 -1973 1369 -1962
rect -45 -2049 349 -2002
rect 1441 -1984 1578 -1950
rect 2689 -1948 2693 -1662
rect 2863 -1718 2894 -1609
rect 2863 -1749 2975 -1718
rect 2944 -1937 2975 -1749
rect 2689 -1952 2827 -1948
rect 2900 -1968 2975 -1937
rect 3459 -1831 4915 -1798
rect 1441 -2038 1475 -1984
rect 3459 -2155 3492 -1831
rect 4882 -1932 4915 -1831
rect 5667 -1932 5704 888
rect 4880 -1969 5704 -1932
rect -435 -2665 -431 -2487
rect -2870 -2669 -431 -2665
rect -2855 -3061 -2850 -2669
rect 932 -2949 964 -2566
rect -1986 -2981 964 -2949
rect -2855 -3066 -2835 -3061
rect -2840 -3088 -2835 -3066
rect -2840 -3094 -2826 -3088
rect -2832 -6427 -2826 -3094
rect -1986 -4655 -1954 -2981
rect 2519 -3165 2566 -2532
rect -1171 -3212 2566 -3165
rect -1708 -4592 -1704 -4484
rect -1879 -4596 -1704 -4592
rect -1879 -4602 -1875 -4596
rect -1287 -4667 -1283 -4493
rect -1171 -4664 -1124 -3212
rect 3990 -3409 4024 -2496
rect 378 -3443 4024 -3409
rect 378 -4121 412 -3443
rect 4280 -3560 4311 -2518
rect 286 -4155 412 -4121
rect 1754 -3591 4311 -3560
rect -145 -4275 201 -4271
rect 197 -4562 201 -4275
rect 197 -4566 215 -4562
rect 211 -4610 215 -4566
rect 286 -4645 320 -4155
rect 963 -4268 1440 -4265
rect -1287 -4671 -1240 -4667
rect 963 -4770 966 -4268
rect 1437 -4315 1440 -4268
rect 1529 -4346 1677 -4342
rect 1673 -4561 1677 -4346
rect 1673 -4565 1686 -4561
rect 1754 -4605 1785 -3591
rect 4581 -3998 4614 -3978
rect 2342 -4030 4614 -3998
rect 2342 -4783 2374 -4030
rect 4581 -4046 4614 -4030
rect 4882 -4046 4915 -1969
rect 4581 -4079 4915 -4046
rect -923 -6427 -917 -5093
rect -2832 -6433 -917 -6427
use and  and_13
timestamp 1669644024
transform 1 0 -1467 0 1 -4544
box -39 -36 185 82
use and  and_12
timestamp 1669644024
transform 1 0 -1889 0 1 -4535
box -39 -36 185 82
use 4bitadder  4bitadder_2
timestamp 1669642337
transform 1 0 -1682 0 1 -5066
box -280 -250 4850 505
use and  and_15
timestamp 1669644024
transform 1 0 1352 0 1 -4393
box -39 -36 185 82
use and  and_14
timestamp 1669644024
transform 1 0 -326 0 1 -4322
box -39 -36 185 82
use 4bitadder  4bitadder_1
timestamp 1669642337
transform 1 0 -538 0 1 -2444
box -280 -250 4850 505
use and  and_11
timestamp 1669644024
transform 1 0 1939 0 1 -1657
box -39 -36 185 82
use and  and_10
timestamp 1669644024
transform 1 0 745 0 1 -1745
box -39 -36 185 82
use and  and_9
timestamp 1669644024
transform 1 0 -129 0 1 -1935
box -39 -36 185 82
use and  and_8
timestamp 1669644024
transform 1 0 -555 0 1 -1642
box -39 -36 185 82
use 4bitadder  4bitadder_0
timestamp 1669642337
transform 1 0 280 0 1 251
box -280 -250 4850 505
use and  and_7
timestamp 1669644024
transform 1 0 3734 0 1 834
box -39 -36 185 82
use and  and_6
timestamp 1669644024
transform 1 0 3444 0 1 830
box -39 -36 185 82
use and  and_5
timestamp 1669644024
transform 1 0 2280 0 1 810
box -39 -36 185 82
use and  and_4
timestamp 1669644024
transform 1 0 1974 0 1 809
box -39 -36 185 82
use and  and_3
timestamp 1669644024
transform 1 0 827 0 1 812
box -39 -36 185 82
use and  and_2
timestamp 1669644024
transform 1 0 555 0 1 810
box -39 -36 185 82
use and  and_1
timestamp 1669644024
transform 1 0 185 0 1 811
box -39 -36 185 82
use and  and_0
timestamp 1669644024
transform 1 0 -135 0 1 812
box -39 -36 185 82
<< labels >>
rlabel space -168 807 -168 807 1 a1_4bitmultiplier
rlabel space -161 781 -161 781 1 b0_4bitmultiplier
rlabel space 153 807 153 807 1 a0_4bitmultiplier
rlabel space 162 778 162 778 1 b1_4bitmultiplier
rlabel space 518 807 518 807 1 a1_4bitmultiplier
rlabel space 531 784 531 784 1 b1_4bitmultiplier
rlabel space 795 808 795 808 1 a2_4bitmultiplier
rlabel space 800 779 800 779 1 b0_4bitmultiplier
rlabel space 1941 805 1941 805 1 a2_4bitmultiplier
rlabel space 1948 778 1948 778 1 b1_4bitmultiplier
rlabel space 2244 805 2244 805 1 a3_4bitmultiplier
rlabel space 2253 780 2253 780 1 b0_4bitmultiplier
rlabel space 3414 824 3414 825 1 a3_4bitmultiplier
rlabel space 3419 797 3419 798 1 b1_4bitmultiplier
rlabel space 470 544 470 544 1 vdd
rlabel space 284 795 284 795 1 gnd
rlabel space 628 794 628 794 1 gnd
rlabel space 940 795 940 795 1 gnd
rlabel space 2069 792 2069 792 1 gnd
rlabel space 2375 793 2375 793 1 gnd
rlabel space 3530 814 3530 814 1 gnd
rlabel space 3833 818 3833 818 1 gnd
rlabel space -587 -1646 -587 -1646 1 a0_4bitmultiplier
rlabel space -581 -1673 -581 -1673 1 b2_4bitmultiplier
rlabel space -162 -1940 -162 -1940 1 a1_4bitmultiplier
rlabel space -156 -1963 -156 -1963 1 b2_4bitmultiplier
rlabel space 712 -1746 712 -1746 1 a2_4bitmultiplier
rlabel space 719 -1774 719 -1774 1 b2_4bitmultiplier
rlabel space 1903 -1663 1903 -1663 1 a3_4bitmultiplier
rlabel space 1914 -1689 1914 -1689 1 b2_4bitmultiplier
rlabel space -1924 -4544 -1924 -4544 1 a0_4bitmultiplier
rlabel space -1916 -4558 -1916 -4558 1 b3_4bitmultiplier
rlabel space -1503 -4550 -1503 -4550 1 a1_4bitmultiplier
rlabel space -1492 -4576 -1492 -4576 1 b3_4bitmultiplier
rlabel space -362 -4328 -362 -4328 1 a2_4bitmultiplier
rlabel space -349 -4353 -349 -4353 1 b3_4bitmultiplier
rlabel space 1321 -4402 1322 -4402 1 a3_4bitmultiplier
rlabel space 1327 -4426 1328 -4426 1 b3_4bitmultiplier
rlabel space -231 -4242 -231 -4242 1 vdd
rlabel space -249 -4339 -249 -4339 1 gnd
rlabel space 640 106 640 106 1 p1_4bitmultiplier
rlabel space -185 -2631 -185 -2631 1 p2_4bitmultiplier
rlabel space -1326 -5225 -1326 -5225 1 p3_4bitmultiplier
rlabel space -197 -5181 -197 -5181 1 p4_4bitmultiplier
rlabel space 1402 -5170 1402 -5170 1 p5_4bitmultiplier
rlabel space 2859 -5128 2859 -5128 1 p6_4bitmultiplier
rlabel space 3146 -5121 3146 -5121 1 p7_4bitmultiplier
<< end >>
