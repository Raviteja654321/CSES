magic
tech scmos
timestamp 1669640031
<< polysilicon >>
rect -24 18 14 21
rect -24 3 -21 18
rect -24 -7 -21 -2
rect 36 -9 38 11
rect -14 -11 38 -9
rect -14 -24 -12 -11
rect -24 -27 -16 -25
<< metal1 >>
rect 40 78 125 82
rect 40 51 44 78
rect 86 49 119 50
rect 85 47 119 49
rect 154 47 185 51
rect 85 46 97 47
rect 85 26 89 46
rect 39 22 89 26
rect 126 19 141 23
rect -39 -2 -24 3
rect -39 -12 -20 -2
rect 10 -15 14 5
rect 137 -15 141 19
rect 10 -19 141 -15
rect -31 -24 -12 -21
rect -31 -29 -16 -24
rect -31 -36 -12 -29
<< metal2 >>
rect 137 47 150 51
<< polycontact >>
rect 119 47 126 51
rect -24 -2 -20 3
rect -16 -29 -12 -24
<< m2contact >>
rect 133 47 137 51
rect 150 47 154 51
use inverter  inverter_0
timestamp 1669639545
transform 1 0 127 0 1 54
box -13 -34 15 28
use nand  nand_0
timestamp 1669639994
transform 1 0 0 0 1 26
box 0 -25 50 29
<< labels >>
rlabel metal1 157 49 157 49 7 v_out_and
rlabel metal1 68 -17 68 -17 1 gnd
rlabel metal1 75 79 75 79 5 vdd
rlabel metal1 -32 -5 -32 -5 1 v_a_and
rlabel metal1 -27 -29 -27 -29 1 v_b_and
<< end >>
