* SPICE3 file created from inverter.ext - technology: scmos

.option scale=1u

M1000 v_out_inv v_in_inv vdd w_n13_n2# pfet w=8 l=2
+  ad=48 pd=28 as=48 ps=28
M1001 v_out_inv v_in_inv gnd Gnd nfet w=8 l=2
+  ad=48 pd=28 as=48 ps=28
C0 w_n13_n2# v_in_inv 3.18fF
C1 gnd Gnd 5.83fF
C2 vdd Gnd 4.70fF
C3 v_in_inv Gnd 5.24fF
