magic
tech scmos
timestamp 1669640721
<< polysilicon >>
rect 25 72 157 74
rect -20 70 15 72
rect -20 31 -18 70
rect -26 29 -18 31
rect -19 24 2 25
rect -26 23 2 24
rect 13 23 15 70
rect 25 51 27 72
rect 61 60 132 62
rect 61 52 63 60
rect 130 52 132 60
rect 155 52 157 72
rect 181 68 232 70
rect 181 31 183 68
rect 230 52 232 68
rect 45 26 62 29
rect 179 30 183 31
rect 102 27 109 30
rect -26 22 -17 23
rect -19 -3 -17 22
rect 13 21 27 23
rect 85 12 89 14
rect 85 -3 87 12
rect 106 -2 109 27
rect 205 1 207 14
rect 203 -1 207 1
rect 268 2 270 16
rect 294 2 296 16
rect 268 0 296 2
rect 203 -2 206 -1
rect -19 -5 89 -3
rect 106 -5 206 -2
rect 268 -16 270 0
<< metal1 >>
rect 305 72 328 78
rect -1 56 4 66
rect 35 55 125 59
rect 165 55 201 59
rect 239 55 265 59
rect 322 43 328 72
rect 322 37 337 43
rect 29 26 39 30
rect 90 27 97 30
rect 161 26 179 30
rect 28 17 32 24
rect 235 23 238 28
rect 244 23 245 28
rect 297 25 335 29
rect 28 13 42 17
rect 1 5 261 9
rect 260 -16 274 -15
rect 260 -20 268 -16
<< metal2 >>
rect 247 72 299 78
rect 305 72 306 78
rect 247 28 255 72
rect 244 23 255 28
rect 42 17 46 18
rect 42 -16 46 13
rect 42 -20 253 -16
rect 268 -20 274 -16
<< polycontact >>
rect 39 26 45 33
rect 97 27 102 31
rect 179 22 184 30
rect 268 -21 274 -16
<< m2contact >>
rect 299 72 305 78
rect 238 23 244 28
rect 42 13 46 17
rect 253 -20 260 -15
use nand  nand_0
timestamp 1669639994
transform 1 0 -11 0 1 30
box 0 -25 50 29
use nand  nand_1
timestamp 1669639994
transform 1 0 50 0 1 30
box 0 -25 50 29
use nand  nand_2
timestamp 1669639994
transform 1 0 119 0 1 30
box 0 -25 50 29
use nand  nand_3
timestamp 1669639994
transform 1 0 194 0 1 30
box 0 -25 50 29
use nand  nand_4
timestamp 1669639994
transform 1 0 257 0 1 31
box 0 -25 50 29
<< labels >>
rlabel metal1 2 62 2 62 5 vdd
rlabel metal1 3 6 3 6 1 gnd
rlabel metal1 331 40 331 40 1 sum_halfadder
rlabel metal1 330 27 330 27 1 carry_halfadder
rlabel polysilicon -24 23 -24 23 3 v_a_halfadder
rlabel polysilicon -24 30 -24 30 3 v_b_halfadder
<< end >>
