magic
tech scmos
timestamp 1669639545
<< nwell >>
rect -13 -2 15 18
<< polysilicon >>
rect -1 12 1 22
rect -1 -4 1 4
rect -3 -7 1 -4
rect -1 -10 1 -7
rect -1 -23 1 -18
<< ndiffusion >>
rect -3 -14 -1 -10
rect -7 -18 -1 -14
rect 1 -14 2 -10
rect 6 -14 7 -10
rect 1 -18 7 -14
<< pdiffusion >>
rect -7 8 -1 12
rect -3 4 -1 8
rect 1 8 7 12
rect 1 4 2 8
rect 6 4 7 8
<< metal1 >>
rect -9 24 10 28
rect -7 8 -3 24
rect 2 -3 6 4
rect 2 -7 8 -3
rect 2 -10 6 -7
rect -7 -30 -3 -14
rect 2 -16 6 -14
rect -9 -34 10 -30
<< ntransistor >>
rect -1 -18 1 -10
<< ptransistor >>
rect -1 4 1 12
<< ndcontact >>
rect -7 -14 -3 -10
rect 2 -14 6 -10
<< pdcontact >>
rect -7 4 -3 8
rect 2 4 6 8
<< labels >>
rlabel metal1 -4 26 -4 26 5 vdd
rlabel metal1 0 -32 0 -32 1 gnd
rlabel polysilicon -2 -6 -2 -6 1 v_in_inv
rlabel metal1 6 -5 6 -5 1 v_out_inv
<< end >>
