* SPICE3 file created from halfadder.ext - technology: scmos

.option scale=1u

M1000 nand_3/a_13_n14# nand_3/v_a_nand gnd Gnd nfet w=4 l=2
+  ad=40 pd=36 as=100 ps=90
M1001 sum_halfadder nand_3/v_b_nand nand_3/a_13_n14# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1002 sum_halfadder nand_3/v_a_nand vdd nand_3/w_0_3# pfet w=8 l=2
+  ad=80 pd=52 as=400 ps=260
M1003 sum_halfadder nand_3/v_b_nand vdd nand_3/w_0_3# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 nand_4/a_13_n14# nand_4/v_b_nand gnd Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1005 carry_halfadder nand_4/v_b_nand nand_4/a_13_n14# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1006 carry_halfadder nand_4/v_b_nand vdd nand_4/w_0_3# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1007 carry_halfadder nand_4/v_b_nand vdd nand_4/w_0_3# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1008 nand_0/a_13_n14# v_a_halfadder gnd Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1009 nand_4/v_b_nand v_b_halfadder nand_0/a_13_n14# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1010 nand_4/v_b_nand v_a_halfadder vdd nand_0/w_0_3# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1011 nand_4/v_b_nand v_b_halfadder vdd nand_0/w_0_3# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1012 nand_1/a_13_n14# nand_4/v_b_nand gnd Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1013 nand_3/v_a_nand v_a_halfadder nand_1/a_13_n14# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1014 nand_3/v_a_nand nand_4/v_b_nand vdd nand_1/w_0_3# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1015 nand_3/v_a_nand v_a_halfadder vdd nand_1/w_0_3# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1016 nand_2/a_13_n14# nand_4/v_b_nand gnd Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1017 nand_3/v_b_nand v_b_halfadder nand_2/a_13_n14# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1018 nand_3/v_b_nand nand_4/v_b_nand vdd nand_2/w_0_3# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1019 nand_3/v_b_nand v_b_halfadder vdd nand_2/w_0_3# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
C0 nand_4/w_0_3# nand_4/v_b_nand 4.92fF
C1 nand_3/v_b_nand nand_3/w_0_3# 2.46fF
C2 nand_1/w_0_3# vdd 2.26fF
C3 nand_1/w_0_3# v_a_halfadder 2.46fF
C4 nand_2/w_0_3# v_b_halfadder 2.46fF
C5 vdd nand_3/w_0_3# 2.26fF
C6 nand_2/w_0_3# vdd 2.26fF
C7 v_b_halfadder nand_0/w_0_3# 6.51fF
C8 nand_0/w_0_3# vdd 2.26fF
C9 nand_0/w_0_3# v_a_halfadder 2.46fF
C10 vdd nand_4/w_0_3# 2.26fF
C11 nand_3/v_a_nand nand_3/w_0_3# 2.46fF
C12 nand_1/w_0_3# nand_4/v_b_nand 2.46fF
C13 nand_2/w_0_3# nand_4/v_b_nand 2.46fF
C14 nand_4/v_b_nand Gnd 106.15fF
C15 v_b_halfadder Gnd 61.26fF
C16 nand_2/a_13_n14# Gnd 2.44fF
C17 nand_3/v_b_nand Gnd 43.65fF
C18 nand_1/a_13_n14# Gnd 2.44fF
C19 gnd Gnd 40.23fF
C20 nand_3/v_a_nand Gnd 27.54fF
C21 nand_0/a_13_n14# Gnd 2.44fF
C22 v_a_halfadder Gnd 54.67fF
C23 nand_4/a_13_n14# Gnd 2.44fF
C24 carry_halfadder Gnd 13.07fF
C25 vdd Gnd 85.63fF
C26 nand_3/a_13_n14# Gnd 2.44fF
C27 sum_halfadder Gnd 20.15fF
