magic
tech scmos
timestamp 1669642337
<< metal1 >>
rect -280 -90 -273 469
rect -198 -48 -190 471
rect 343 381 358 404
rect 343 352 358 355
rect 428 372 460 413
rect 490 373 522 425
rect 1889 397 1909 477
rect 428 351 429 372
rect 516 363 522 373
rect 1476 342 1489 389
rect 1487 328 1489 342
rect 1982 383 2002 480
rect 3352 436 3388 505
rect 1889 327 1909 341
rect 3075 344 3087 388
rect 3352 368 3353 436
rect 3385 368 3388 436
rect 3352 365 3388 368
rect 3431 426 3467 498
rect 3463 358 3467 426
rect 3083 325 3087 344
rect 4536 357 4549 401
rect 4546 340 4549 357
rect 1520 298 2201 303
rect 52 292 607 296
rect 2196 292 2201 298
rect 3120 297 3659 302
rect 3654 295 3659 297
rect 42 233 46 241
rect 52 233 56 292
rect 3654 290 3666 295
rect 383 243 554 246
rect 2034 245 2150 249
rect 42 229 56 233
rect 381 239 554 243
rect 42 77 46 229
rect -110 54 -81 55
rect -110 50 -1 54
rect 381 51 387 239
rect 2035 152 2039 245
rect 3523 244 3613 248
rect 3523 243 3605 244
rect 3609 243 3613 244
rect 3523 239 3613 243
rect 3523 155 3527 239
rect 1777 148 2039 152
rect 3375 151 3527 155
rect 454 77 536 85
rect 355 47 387 51
rect -7 46 0 47
rect -87 45 0 46
rect -89 44 0 45
rect -80 43 0 44
rect -80 42 5 43
rect -80 41 -2 42
rect -110 -48 -102 23
rect -198 -56 -102 -48
rect -89 -90 -82 24
rect 39 -43 43 31
rect 442 3 450 69
rect 448 -11 450 3
rect 442 -13 450 -11
rect 490 29 494 44
rect 512 36 539 44
rect 490 3 498 29
rect 497 -11 498 3
rect 490 -12 498 -11
rect 615 -43 619 -29
rect 1549 -33 1556 84
rect 1914 80 2133 88
rect 3323 78 3353 86
rect 1900 10 1908 63
rect 3323 56 3331 78
rect 3386 78 3593 86
rect 1997 39 2136 47
rect 1972 12 1980 35
rect 3401 37 3440 45
rect 3473 37 3596 45
rect 3277 -3 3284 2
rect 3663 -3 3670 5
rect 2900 -10 3670 -3
rect 3663 -11 3670 -10
rect 1972 -14 1980 -11
rect 4528 -13 4562 -10
rect 2204 -33 2216 -22
rect 1549 -40 2216 -33
rect 4528 -34 4536 -13
rect 4545 -34 4562 -13
rect 39 -47 619 -43
rect 2204 -44 2211 -40
rect 3307 -51 3357 -50
rect 3307 -54 3320 -51
rect 1470 -56 1493 -55
rect 346 -58 364 -57
rect 346 -63 348 -58
rect 362 -63 364 -58
rect 346 -72 364 -63
rect 1470 -67 1478 -56
rect 1487 -60 1493 -56
rect 1487 -67 1502 -60
rect -280 -97 -82 -90
rect 345 -250 367 -72
rect 441 -74 452 -69
rect 441 -88 443 -74
rect 450 -88 452 -74
rect 441 -93 452 -88
rect 487 -84 491 -70
rect 487 -93 498 -84
rect 423 -146 461 -93
rect 484 -146 522 -93
rect 1470 -163 1502 -67
rect 1880 -77 1916 -72
rect 1880 -100 1898 -77
rect 1912 -100 1916 -77
rect 1880 -155 1916 -100
rect 1958 -82 1994 -72
rect 1958 -105 1969 -82
rect 1983 -105 1994 -82
rect 1958 -155 1994 -105
rect 3057 -78 3072 -56
rect 3086 -78 3104 -56
rect 3057 -135 3104 -78
rect 3308 -76 3320 -54
rect 3341 -76 3357 -51
rect 3308 -138 3357 -76
rect 3372 -76 3377 -52
rect 3398 -76 3416 -52
rect 3372 -111 3416 -76
rect 4528 -100 4562 -34
rect 4818 -18 4849 -4
rect 4818 -23 4820 -18
rect 4836 -23 4849 -18
rect 4818 -86 4849 -23
rect 4818 -99 4850 -86
rect 3370 -139 3417 -111
rect 4818 -113 4849 -99
rect 3372 -140 3409 -139
<< metal2 >>
rect 345 381 358 384
rect 436 372 456 375
rect 491 373 511 399
rect 345 100 358 355
rect 345 87 358 88
rect 436 87 456 344
rect 454 69 456 87
rect 347 65 362 67
rect 436 66 456 69
rect 347 60 349 65
rect -115 45 -110 50
rect -100 45 -97 50
rect -115 28 -97 45
rect -115 23 -110 28
rect -100 23 -97 28
rect -91 39 -90 44
rect -80 39 -77 44
rect -91 29 -77 39
rect -91 24 -90 29
rect -80 24 -77 29
rect 347 -58 362 60
rect 491 47 511 345
rect 1477 342 1488 344
rect 1487 328 1488 342
rect 1477 257 1488 328
rect 1477 251 1478 257
rect 1487 251 1488 257
rect 593 241 597 246
rect 1477 245 1488 251
rect 1887 341 1888 397
rect 491 29 494 47
rect 491 25 511 29
rect 442 3 450 4
rect 448 -11 450 3
rect 347 -63 348 -58
rect 347 -65 362 -63
rect 442 -74 450 -11
rect 442 -88 443 -74
rect 489 3 498 8
rect 489 -11 490 3
rect 497 -11 498 3
rect 489 -70 498 -11
rect 489 -84 491 -70
rect 1478 -56 1486 245
rect 1887 119 1911 341
rect 1974 327 1978 364
rect 3436 426 3466 432
rect 3385 368 3386 410
rect 1887 68 1890 119
rect 1974 55 1998 327
rect 1997 35 1998 55
rect 3074 325 3075 344
rect 3074 260 3083 325
rect 3074 253 3075 260
rect 1898 10 1911 11
rect 1478 -76 1486 -67
rect 489 -86 498 -84
rect 1898 -77 1911 -13
rect 442 -89 450 -88
rect 1968 -82 1981 -11
rect 3074 -55 3083 253
rect 3356 92 3386 368
rect 3463 369 3466 426
rect 3463 358 3468 369
rect 3436 99 3468 358
rect 4546 340 4547 357
rect 4536 259 4547 340
rect 4536 251 4537 259
rect 4546 251 4547 259
rect 4536 248 4547 251
rect 3341 28 3342 56
rect 3319 -51 3342 28
rect 3319 -75 3320 -51
rect 3341 -75 3342 -51
rect 3374 52 3397 58
rect 3374 24 3375 52
rect 3438 51 3468 99
rect 3438 36 3440 51
rect 3374 -51 3397 24
rect 4537 -13 4545 248
rect 4820 149 4821 154
rect 4820 -18 4837 149
rect 4836 -23 4837 -18
rect 4820 -25 4837 -23
rect 4537 -35 4545 -34
rect 3374 -73 3377 -51
rect 3074 -79 3083 -78
rect 1898 -111 1911 -100
rect 1968 -105 1969 -82
rect 1968 -112 1981 -105
<< polycontact >>
rect -1 50 5 54
rect 0 43 6 47
<< m2contact >>
rect 342 355 358 381
rect 429 344 461 372
rect 484 345 516 373
rect 1476 328 1487 342
rect 1888 341 1912 397
rect 1978 327 2002 383
rect 3353 368 3385 436
rect 3431 358 3463 426
rect 3075 325 3083 344
rect 4536 340 4546 357
rect 1478 251 1487 257
rect 3075 253 3083 260
rect 4537 251 4546 259
rect 345 88 359 100
rect 349 60 363 65
rect 4821 149 4837 154
rect 436 69 454 87
rect -110 45 -100 50
rect -90 39 -80 44
rect -110 23 -100 28
rect -90 24 -80 29
rect 441 -11 448 3
rect 494 29 512 47
rect 490 -11 497 3
rect 1890 63 1914 119
rect 3353 75 3386 92
rect 1971 35 1997 55
rect 3315 28 3341 56
rect 3375 24 3401 52
rect 3440 34 3473 51
rect 1898 -13 1912 10
rect 1968 -11 1982 12
rect 4536 -34 4545 -13
rect 348 -63 362 -58
rect 1478 -67 1487 -56
rect 443 -88 450 -74
rect 491 -84 498 -70
rect 1898 -100 1912 -77
rect 1969 -105 1983 -82
rect 3072 -78 3086 -55
rect 3320 -76 3341 -51
rect 3377 -76 3398 -51
rect 4820 -23 4836 -18
use fulladder  fulladder_2
timestamp 1669640721
transform 1 0 3640 0 1 14
box -55 -48 1200 290
use fulladder  fulladder_1
timestamp 1669640721
transform 1 0 2180 0 1 16
box -55 -48 1200 290
use fulladder  fulladder_0
timestamp 1669640721
transform 1 0 583 0 1 13
box -55 -48 1200 290
use halfadder  halfadder_0
timestamp 1669640721
transform 1 0 25 0 1 22
box -26 -21 337 78
<< labels >>
rlabel metal1 56 294 56 294 1 vdd
rlabel metal1 2031 300 2031 300 1 vdd
rlabel metal1 3442 298 3442 298 1 vdd
rlabel metal1 308 -46 308 -46 1 gnd
rlabel metal1 1870 -37 1870 -37 1 gnd
rlabel metal1 3282 -9 3282 -6 1 gnd
rlabel metal1 350 -76 350 -76 1 s0_4bitadder
rlabel metal1 446 -103 446 -103 1 a1_4bitadder
rlabel metal1 493 -103 493 -103 1 b1_4bitadder
rlabel metal1 354 -211 354 -211 1 s0_4bitadder
rlabel metal1 1484 -143 1484 -142 1 s1_4bitadder
rlabel metal1 3068 -113 3068 -113 1 s2_4bitadder
rlabel metal1 1981 -132 1981 -132 1 b2_4bitadder
rlabel metal1 1896 -125 1896 -125 1 a2_4bitadder
rlabel metal1 3325 -107 3325 -107 1 a3_4bitadder
rlabel metal1 3385 -112 3385 -112 1 b3_4bitadder
rlabel metal1 4543 -78 4543 -78 1 s3_4bitadder
rlabel metal1 4833 -73 4833 -73 1 c_4bitadder
rlabel metal1 -108 12 -108 12 1 a0_4bitadder
rlabel metal1 -86 13 -86 13 1 b0_4bitadder
rlabel metal1 351 398 351 398 1 s0_4bitadder
rlabel metal1 1479 374 1479 374 1 s1_4bitadder
rlabel metal1 3078 366 3078 366 1 s2_4bitadder
rlabel metal1 4542 376 4542 376 1 s3_4bitadder
rlabel metal1 3371 480 3371 480 1 a3_4bitadder
rlabel metal1 3452 457 3452 457 1 b3_4bitadder
rlabel metal1 1898 432 1898 432 1 a2_4bitadder
rlabel metal1 1898 432 1898 432 1 b2_4bitadder
rlabel metal1 446 391 448 392 1 a1_4bitadder
rlabel metal1 446 391 448 392 1 b1_4bitadder
rlabel metal1 511 406 511 406 1 b1_4bitadder
rlabel metal1 -277 452 -276 453 3 b0_4bitadder
rlabel metal1 -194 453 -194 453 1 a0_4bitadder
rlabel metal1 1992 421 1992 421 1 b2_4bitadder
<< end >>
