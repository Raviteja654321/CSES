magic
tech scmos
timestamp 1669639994
<< nwell >>
rect 0 3 49 20
<< polysilicon >>
rect 11 14 13 24
rect 36 14 38 24
rect 11 -10 13 6
rect 36 -10 38 6
rect 11 -18 13 -14
rect 36 -18 38 -14
<< ndiffusion >>
rect 10 -14 11 -10
rect 13 -14 14 -10
rect 35 -14 36 -10
rect 38 -14 39 -10
<< pdiffusion >>
rect 10 6 11 14
rect 13 6 14 14
rect 35 6 36 14
rect 38 6 39 14
<< metal1 >>
rect 1 25 50 29
rect 6 14 10 25
rect 31 14 35 25
rect 14 1 18 6
rect 39 1 43 6
rect 14 -3 43 1
rect 39 -10 43 -3
rect 18 -14 31 -10
rect 6 -21 10 -14
rect 0 -25 16 -21
<< ntransistor >>
rect 11 -14 13 -10
rect 36 -14 38 -10
<< ptransistor >>
rect 11 6 13 14
rect 36 6 38 14
<< ndcontact >>
rect 6 -14 10 -10
rect 14 -14 18 -10
rect 31 -14 35 -10
rect 39 -14 43 -10
<< pdcontact >>
rect 6 6 10 14
rect 14 6 18 14
rect 31 6 35 14
rect 39 6 43 14
<< labels >>
rlabel metal1 23 27 23 27 5 vdd
rlabel metal1 9 -23 9 -23 1 gnd
rlabel metal1 41 -2 41 -2 1 v_out_nand
<< end >>
