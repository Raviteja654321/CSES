magic
tech scmos
timestamp 1669640721
<< polysilicon >>
rect 499 228 500 232
rect 505 228 508 232
rect 499 223 505 225
rect 499 209 501 223
rect 496 207 501 209
rect -43 68 -42 70
rect -35 68 -14 70
rect -16 53 -14 68
rect -16 51 -5 53
rect -16 44 -5 46
rect -42 28 -39 30
rect -16 30 -14 44
rect -32 28 -14 30
<< metal1 >>
rect 528 285 945 290
rect 528 284 533 285
rect 17 279 533 284
rect -38 229 -1 233
rect 9 229 14 233
rect -38 228 14 229
rect 17 122 22 279
rect 528 262 533 279
rect 890 238 910 244
rect 74 227 75 233
rect 85 232 508 233
rect 85 228 500 232
rect 505 228 508 232
rect 85 227 508 228
rect 860 226 889 230
rect 484 211 498 212
rect 456 209 498 211
rect 456 205 492 209
rect 496 205 498 209
rect 17 117 23 122
rect 17 112 25 117
rect 18 83 23 112
rect -55 65 -42 72
rect 456 65 462 205
rect 484 203 498 205
rect 544 173 548 210
rect 544 141 553 173
rect 552 131 553 141
rect 885 132 889 226
rect 940 187 945 285
rect 1161 135 1200 139
rect 885 128 910 132
rect 915 128 918 132
rect 899 123 917 125
rect 899 119 910 123
rect 915 119 917 123
rect 899 117 917 119
rect 899 114 903 117
rect -55 64 -35 65
rect 349 59 462 65
rect 477 110 903 114
rect 477 51 481 110
rect 997 71 1011 97
rect 551 64 1011 71
rect 350 47 481 51
rect -52 25 -39 31
rect -52 23 -32 25
rect 26 -40 30 31
rect 722 -40 729 64
rect 25 -46 729 -40
rect 722 -48 729 -46
<< metal2 >>
rect 866 238 882 244
rect 9 233 86 234
rect 9 229 75 233
rect -1 227 75 229
rect 85 227 86 233
rect 1124 135 1150 139
rect 1161 135 1163 139
rect 544 73 551 130
<< polycontact >>
rect 500 228 505 232
rect 492 205 496 209
rect 910 128 915 132
rect 910 119 915 123
rect -42 65 -35 72
rect -39 25 -32 31
<< m2contact >>
rect -1 229 9 235
rect 858 238 866 244
rect 882 238 890 244
rect 75 227 85 233
rect 542 130 552 141
rect 1113 135 1124 139
rect 1150 135 1161 139
rect 541 62 551 73
use or  or_0
timestamp 1669631468
transform 1 0 976 0 1 140
box -66 -52 147 53
use halfadder  halfadder_0
timestamp 1669640721
transform 1 0 19 0 1 22
box -26 -21 337 78
use halfadder  halfadder_1
timestamp 1669640721
transform 1 0 529 0 1 201
box -26 -21 337 78
<< labels >>
rlabel polycontact -38 29 -38 29 3 v_b_fulladder
rlabel polycontact -40 69 -40 69 3 v_a_fulladder
rlabel metal1 906 241 906 241 1 sum_fulladder
rlabel metal1 1186 137 1186 137 1 carry_fulladder
rlabel metal1 480 229 480 229 1 c_in_fulladder
rlabel space 574 258 574 258 1 vdd
rlabel metal1 530 286 530 286 5 vdd
rlabel metal1 545 172 545 172 1 gnd
rlabel metal1 21 110 21 110 1 vdd
rlabel metal1 27 -9 27 -9 1 gnd
rlabel space 929 178 929 178 1 vdd
rlabel metal1 1006 94 1006 94 1 gnd
rlabel metal1 -31 231 -31 231 1 c_in_fulladder
rlabel metal1 18 281 18 281 1 vdd
rlabel metal1 345 -43 345 -43 1 gnd
<< end >>
