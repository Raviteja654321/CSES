* SPICE3 file created from 4bitadder.ext - technology: scmos

.option scale=1u

M1000 halfadder_0/nand_3/a_13_n14# halfadder_0/nand_1/v_out_nand gnd Gnd nfet w=4 l=2
+  ad=40 pd=36 as=1372 ps=978
M1001 s0_4bitadder halfadder_0/nand_2/v_out_nand halfadder_0/nand_3/a_13_n14# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1002 s0_4bitadder halfadder_0/nand_1/v_out_nand vdd halfadder_0/nand_3/w_0_3# pfet w=8 l=2
+  ad=80 pd=52 as=3259 ps=2060
M1003 s0_4bitadder halfadder_0/nand_2/v_out_nand vdd halfadder_0/nand_3/w_0_3# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 halfadder_0/nand_4/a_13_n14# halfadder_0/nand_0/v_out_nand gnd Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1005 fulladder_0/c_in_fulladder halfadder_0/nand_0/v_out_nand halfadder_0/nand_4/a_13_n14# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1006 fulladder_0/c_in_fulladder halfadder_0/nand_0/v_out_nand vdd halfadder_0/nand_4/w_0_3# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1007 fulladder_0/c_in_fulladder halfadder_0/nand_0/v_out_nand vdd halfadder_0/nand_4/w_0_3# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1008 halfadder_0/nand_0/a_13_n14# b0_4bitadder gnd Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1009 halfadder_0/nand_0/v_out_nand a0_4bitadder halfadder_0/nand_0/a_13_n14# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1010 halfadder_0/nand_0/v_out_nand b0_4bitadder vdd halfadder_0/nand_0/w_0_3# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1011 halfadder_0/nand_0/v_out_nand a0_4bitadder vdd halfadder_0/nand_0/w_0_3# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1012 halfadder_0/nand_1/a_13_n14# halfadder_0/nand_0/v_out_nand gnd Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1013 halfadder_0/nand_1/v_out_nand b0_4bitadder halfadder_0/nand_1/a_13_n14# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1014 halfadder_0/nand_1/v_out_nand halfadder_0/nand_0/v_out_nand vdd halfadder_0/nand_1/w_0_3# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1015 halfadder_0/nand_1/v_out_nand b0_4bitadder vdd halfadder_0/nand_1/w_0_3# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1016 halfadder_0/nand_2/a_13_n14# halfadder_0/nand_0/v_out_nand gnd Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1017 halfadder_0/nand_2/v_out_nand a0_4bitadder halfadder_0/nand_2/a_13_n14# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1018 halfadder_0/nand_2/v_out_nand halfadder_0/nand_0/v_out_nand vdd halfadder_0/nand_2/w_0_3# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1019 halfadder_0/nand_2/v_out_nand a0_4bitadder vdd halfadder_0/nand_2/w_0_3# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1020 fulladder_0/halfadder_0/nand_3/a_13_n14# fulladder_0/halfadder_0/nand_1/v_out_nand gnd Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1021 fulladder_0/halfadder_1/v_a_halfadder fulladder_0/halfadder_0/nand_2/v_out_nand fulladder_0/halfadder_0/nand_3/a_13_n14# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1022 fulladder_0/halfadder_1/v_a_halfadder fulladder_0/halfadder_0/nand_1/v_out_nand vdd fulladder_0/halfadder_0/nand_3/w_0_3# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1023 fulladder_0/halfadder_1/v_a_halfadder fulladder_0/halfadder_0/nand_2/v_out_nand vdd fulladder_0/halfadder_0/nand_3/w_0_3# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1024 fulladder_0/halfadder_0/nand_4/a_13_n14# fulladder_0/halfadder_0/nand_0/v_out_nand gnd Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1025 fulladder_0/or_0/v_b_or fulladder_0/halfadder_0/nand_0/v_out_nand fulladder_0/halfadder_0/nand_4/a_13_n14# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1026 fulladder_0/or_0/v_b_or fulladder_0/halfadder_0/nand_0/v_out_nand vdd fulladder_0/halfadder_0/nand_4/w_0_3# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1027 fulladder_0/or_0/v_b_or fulladder_0/halfadder_0/nand_0/v_out_nand vdd fulladder_0/halfadder_0/nand_4/w_0_3# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1028 fulladder_0/halfadder_0/nand_0/a_13_n14# b1_4bitadder gnd Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1029 fulladder_0/halfadder_0/nand_0/v_out_nand b1_4bitadder fulladder_0/halfadder_0/nand_0/a_13_n14# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1030 fulladder_0/halfadder_0/nand_0/v_out_nand b1_4bitadder vdd fulladder_0/halfadder_0/nand_0/w_0_3# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1031 fulladder_0/halfadder_0/nand_0/v_out_nand b1_4bitadder vdd fulladder_0/halfadder_0/nand_0/w_0_3# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1032 fulladder_0/halfadder_0/nand_1/a_13_n14# fulladder_0/halfadder_0/nand_0/v_out_nand gnd Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1033 fulladder_0/halfadder_0/nand_1/v_out_nand b1_4bitadder fulladder_0/halfadder_0/nand_1/a_13_n14# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1034 fulladder_0/halfadder_0/nand_1/v_out_nand fulladder_0/halfadder_0/nand_0/v_out_nand vdd fulladder_0/halfadder_0/nand_1/w_0_3# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1035 fulladder_0/halfadder_0/nand_1/v_out_nand b1_4bitadder vdd fulladder_0/halfadder_0/nand_1/w_0_3# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1036 fulladder_0/halfadder_0/nand_2/a_13_n14# fulladder_0/halfadder_0/nand_0/v_out_nand gnd Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1037 fulladder_0/halfadder_0/nand_2/v_out_nand b1_4bitadder fulladder_0/halfadder_0/nand_2/a_13_n14# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1038 fulladder_0/halfadder_0/nand_2/v_out_nand fulladder_0/halfadder_0/nand_0/v_out_nand vdd fulladder_0/halfadder_0/nand_2/w_0_3# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1039 fulladder_0/halfadder_0/nand_2/v_out_nand b1_4bitadder vdd fulladder_0/halfadder_0/nand_2/w_0_3# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1040 fulladder_0/halfadder_1/nand_3/a_13_n14# fulladder_0/halfadder_1/nand_1/v_out_nand gnd Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1041 s1_4bitadder fulladder_0/halfadder_1/nand_2/v_out_nand fulladder_0/halfadder_1/nand_3/a_13_n14# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1042 s1_4bitadder fulladder_0/halfadder_1/nand_1/v_out_nand vdd fulladder_0/halfadder_1/nand_3/w_0_3# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1043 s1_4bitadder fulladder_0/halfadder_1/nand_2/v_out_nand vdd fulladder_0/halfadder_1/nand_3/w_0_3# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1044 fulladder_0/halfadder_1/nand_4/a_13_n14# fulladder_0/halfadder_1/nand_0/v_out_nand gnd Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1045 fulladder_0/or_0/v_a_or fulladder_0/halfadder_1/nand_0/v_out_nand fulladder_0/halfadder_1/nand_4/a_13_n14# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1046 fulladder_0/or_0/v_a_or fulladder_0/halfadder_1/nand_0/v_out_nand vdd fulladder_0/halfadder_1/nand_4/w_0_3# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1047 fulladder_0/or_0/v_a_or fulladder_0/halfadder_1/nand_0/v_out_nand vdd fulladder_0/halfadder_1/nand_4/w_0_3# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1048 fulladder_0/halfadder_1/nand_0/a_13_n14# fulladder_0/halfadder_1/v_a_halfadder gnd Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1049 fulladder_0/halfadder_1/nand_0/v_out_nand fulladder_0/c_in_fulladder fulladder_0/halfadder_1/nand_0/a_13_n14# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1050 fulladder_0/halfadder_1/nand_0/v_out_nand fulladder_0/halfadder_1/v_a_halfadder vdd fulladder_0/halfadder_1/nand_0/w_0_3# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1051 fulladder_0/halfadder_1/nand_0/v_out_nand fulladder_0/c_in_fulladder vdd fulladder_0/halfadder_1/nand_0/w_0_3# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1052 fulladder_0/halfadder_1/nand_1/a_13_n14# fulladder_0/halfadder_1/nand_0/v_out_nand gnd Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1053 fulladder_0/halfadder_1/nand_1/v_out_nand fulladder_0/halfadder_1/v_a_halfadder fulladder_0/halfadder_1/nand_1/a_13_n14# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1054 fulladder_0/halfadder_1/nand_1/v_out_nand fulladder_0/halfadder_1/nand_0/v_out_nand vdd fulladder_0/halfadder_1/nand_1/w_0_3# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1055 fulladder_0/halfadder_1/nand_1/v_out_nand fulladder_0/halfadder_1/v_a_halfadder vdd fulladder_0/halfadder_1/nand_1/w_0_3# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1056 fulladder_0/halfadder_1/nand_2/a_13_n14# fulladder_0/halfadder_1/nand_0/v_out_nand gnd Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1057 fulladder_0/halfadder_1/nand_2/v_out_nand fulladder_0/c_in_fulladder fulladder_0/halfadder_1/nand_2/a_13_n14# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1058 fulladder_0/halfadder_1/nand_2/v_out_nand fulladder_0/halfadder_1/nand_0/v_out_nand vdd fulladder_0/halfadder_1/nand_2/w_0_3# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1059 fulladder_0/halfadder_1/nand_2/v_out_nand fulladder_0/c_in_fulladder vdd fulladder_0/halfadder_1/nand_2/w_0_3# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1060 fulladder_0/or_0/a_n15_n30# fulladder_0/or_0/v_b_or gnd Gnd nfet w=12 l=3
+  ad=156 pd=74 as=0 ps=0
M1061 fulladder_0/or_0/a_n15_n30# fulladder_0/or_0/v_a_or gnd Gnd nfet w=12 l=3
+  ad=0 pd=0 as=0 ps=0
M1062 fulladder_1/c_in_fulladder fulladder_0/or_0/a_n15_n30# gnd Gnd nfet w=16 l=3
+  ad=84 pd=44 as=0 ps=0
M1063 fulladder_0/or_0/a_n15_10# fulladder_0/or_0/v_a_or vdd fulladder_0/or_0/w_n32_2# pfet w=12 l=3
+  ad=156 pd=74 as=0 ps=0
M1064 vdd fulladder_0/or_0/a_n15_n30# fulladder_1/c_in_fulladder fulladder_0/or_0/w_78_2# pfet w=16 l=3
+  ad=0 pd=0 as=80 ps=42
M1065 fulladder_0/or_0/a_n15_n30# fulladder_0/or_0/v_b_or fulladder_0/or_0/a_n15_10# fulladder_0/or_0/w_n32_2# pfet w=12 l=3
+  ad=72 pd=36 as=0 ps=0
M1066 fulladder_1/halfadder_0/nand_3/a_13_n14# fulladder_1/halfadder_0/nand_1/v_out_nand gnd Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1067 fulladder_1/halfadder_1/v_a_halfadder fulladder_1/halfadder_0/nand_2/v_out_nand fulladder_1/halfadder_0/nand_3/a_13_n14# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1068 fulladder_1/halfadder_1/v_a_halfadder fulladder_1/halfadder_0/nand_1/v_out_nand vdd fulladder_1/halfadder_0/nand_3/w_0_3# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1069 fulladder_1/halfadder_1/v_a_halfadder fulladder_1/halfadder_0/nand_2/v_out_nand vdd fulladder_1/halfadder_0/nand_3/w_0_3# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1070 fulladder_1/halfadder_0/nand_4/a_13_n14# fulladder_1/halfadder_0/nand_0/v_out_nand gnd Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1071 fulladder_1/or_0/v_b_or fulladder_1/halfadder_0/nand_0/v_out_nand fulladder_1/halfadder_0/nand_4/a_13_n14# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1072 fulladder_1/or_0/v_b_or fulladder_1/halfadder_0/nand_0/v_out_nand vdd fulladder_1/halfadder_0/nand_4/w_0_3# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1073 fulladder_1/or_0/v_b_or fulladder_1/halfadder_0/nand_0/v_out_nand vdd fulladder_1/halfadder_0/nand_4/w_0_3# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1074 fulladder_1/halfadder_0/nand_0/a_13_n14# b2_4bitadder gnd Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1075 fulladder_1/halfadder_0/nand_0/v_out_nand b2_4bitadder fulladder_1/halfadder_0/nand_0/a_13_n14# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1076 fulladder_1/halfadder_0/nand_0/v_out_nand b2_4bitadder vdd fulladder_1/halfadder_0/nand_0/w_0_3# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1077 fulladder_1/halfadder_0/nand_0/v_out_nand b2_4bitadder vdd fulladder_1/halfadder_0/nand_0/w_0_3# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1078 fulladder_1/halfadder_0/nand_1/a_13_n14# fulladder_1/halfadder_0/nand_0/v_out_nand gnd Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1079 fulladder_1/halfadder_0/nand_1/v_out_nand b2_4bitadder fulladder_1/halfadder_0/nand_1/a_13_n14# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1080 fulladder_1/halfadder_0/nand_1/v_out_nand fulladder_1/halfadder_0/nand_0/v_out_nand vdd fulladder_1/halfadder_0/nand_1/w_0_3# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1081 fulladder_1/halfadder_0/nand_1/v_out_nand b2_4bitadder vdd fulladder_1/halfadder_0/nand_1/w_0_3# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1082 fulladder_1/halfadder_0/nand_2/a_13_n14# fulladder_1/halfadder_0/nand_0/v_out_nand gnd Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1083 fulladder_1/halfadder_0/nand_2/v_out_nand b2_4bitadder fulladder_1/halfadder_0/nand_2/a_13_n14# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1084 fulladder_1/halfadder_0/nand_2/v_out_nand fulladder_1/halfadder_0/nand_0/v_out_nand vdd fulladder_1/halfadder_0/nand_2/w_0_3# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1085 fulladder_1/halfadder_0/nand_2/v_out_nand b2_4bitadder vdd fulladder_1/halfadder_0/nand_2/w_0_3# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1086 fulladder_1/halfadder_1/nand_3/a_13_n14# fulladder_1/halfadder_1/nand_1/v_out_nand gnd Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1087 s2_4bitadder fulladder_1/halfadder_1/nand_2/v_out_nand fulladder_1/halfadder_1/nand_3/a_13_n14# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1088 s2_4bitadder fulladder_1/halfadder_1/nand_1/v_out_nand vdd fulladder_1/halfadder_1/nand_3/w_0_3# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1089 s2_4bitadder fulladder_1/halfadder_1/nand_2/v_out_nand vdd fulladder_1/halfadder_1/nand_3/w_0_3# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1090 fulladder_1/halfadder_1/nand_4/a_13_n14# fulladder_1/halfadder_1/nand_0/v_out_nand gnd Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1091 fulladder_1/or_0/v_a_or fulladder_1/halfadder_1/nand_0/v_out_nand fulladder_1/halfadder_1/nand_4/a_13_n14# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1092 fulladder_1/or_0/v_a_or fulladder_1/halfadder_1/nand_0/v_out_nand vdd fulladder_1/halfadder_1/nand_4/w_0_3# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1093 fulladder_1/or_0/v_a_or fulladder_1/halfadder_1/nand_0/v_out_nand vdd fulladder_1/halfadder_1/nand_4/w_0_3# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1094 fulladder_1/halfadder_1/nand_0/a_13_n14# fulladder_1/halfadder_1/v_a_halfadder gnd Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1095 fulladder_1/halfadder_1/nand_0/v_out_nand fulladder_1/c_in_fulladder fulladder_1/halfadder_1/nand_0/a_13_n14# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1096 fulladder_1/halfadder_1/nand_0/v_out_nand fulladder_1/halfadder_1/v_a_halfadder vdd fulladder_1/halfadder_1/nand_0/w_0_3# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1097 fulladder_1/halfadder_1/nand_0/v_out_nand fulladder_1/c_in_fulladder vdd fulladder_1/halfadder_1/nand_0/w_0_3# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1098 fulladder_1/halfadder_1/nand_1/a_13_n14# fulladder_1/halfadder_1/nand_0/v_out_nand gnd Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1099 fulladder_1/halfadder_1/nand_1/v_out_nand fulladder_1/halfadder_1/v_a_halfadder fulladder_1/halfadder_1/nand_1/a_13_n14# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1100 fulladder_1/halfadder_1/nand_1/v_out_nand fulladder_1/halfadder_1/nand_0/v_out_nand vdd fulladder_1/halfadder_1/nand_1/w_0_3# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1101 fulladder_1/halfadder_1/nand_1/v_out_nand fulladder_1/halfadder_1/v_a_halfadder vdd fulladder_1/halfadder_1/nand_1/w_0_3# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1102 fulladder_1/halfadder_1/nand_2/a_13_n14# fulladder_1/halfadder_1/nand_0/v_out_nand gnd Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1103 fulladder_1/halfadder_1/nand_2/v_out_nand fulladder_1/c_in_fulladder fulladder_1/halfadder_1/nand_2/a_13_n14# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1104 fulladder_1/halfadder_1/nand_2/v_out_nand fulladder_1/halfadder_1/nand_0/v_out_nand vdd fulladder_1/halfadder_1/nand_2/w_0_3# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1105 fulladder_1/halfadder_1/nand_2/v_out_nand fulladder_1/c_in_fulladder vdd fulladder_1/halfadder_1/nand_2/w_0_3# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1106 fulladder_1/or_0/a_n15_n30# fulladder_1/or_0/v_b_or gnd Gnd nfet w=12 l=3
+  ad=156 pd=74 as=0 ps=0
M1107 fulladder_1/or_0/a_n15_n30# fulladder_1/or_0/v_a_or gnd Gnd nfet w=12 l=3
+  ad=0 pd=0 as=0 ps=0
M1108 fulladder_2/c_in_fulladder fulladder_1/or_0/a_n15_n30# gnd Gnd nfet w=16 l=3
+  ad=84 pd=44 as=0 ps=0
M1109 fulladder_1/or_0/a_n15_10# fulladder_1/or_0/v_a_or vdd fulladder_1/or_0/w_n32_2# pfet w=12 l=3
+  ad=156 pd=74 as=0 ps=0
M1110 vdd fulladder_1/or_0/a_n15_n30# fulladder_2/c_in_fulladder fulladder_1/or_0/w_78_2# pfet w=16 l=3
+  ad=0 pd=0 as=80 ps=42
M1111 fulladder_1/or_0/a_n15_n30# fulladder_1/or_0/v_b_or fulladder_1/or_0/a_n15_10# fulladder_1/or_0/w_n32_2# pfet w=12 l=3
+  ad=72 pd=36 as=0 ps=0
M1112 fulladder_2/halfadder_0/nand_3/a_13_n14# fulladder_2/halfadder_0/nand_1/v_out_nand gnd Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1113 fulladder_2/halfadder_1/v_a_halfadder fulladder_2/halfadder_0/nand_2/v_out_nand fulladder_2/halfadder_0/nand_3/a_13_n14# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1114 fulladder_2/halfadder_1/v_a_halfadder fulladder_2/halfadder_0/nand_1/v_out_nand vdd fulladder_2/halfadder_0/nand_3/w_0_3# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1115 fulladder_2/halfadder_1/v_a_halfadder fulladder_2/halfadder_0/nand_2/v_out_nand vdd fulladder_2/halfadder_0/nand_3/w_0_3# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1116 fulladder_2/halfadder_0/nand_4/a_13_n14# fulladder_2/halfadder_0/nand_0/v_out_nand gnd Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1117 fulladder_2/or_0/v_b_or fulladder_2/halfadder_0/nand_0/v_out_nand fulladder_2/halfadder_0/nand_4/a_13_n14# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1118 fulladder_2/or_0/v_b_or fulladder_2/halfadder_0/nand_0/v_out_nand vdd fulladder_2/halfadder_0/nand_4/w_0_3# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1119 fulladder_2/or_0/v_b_or fulladder_2/halfadder_0/nand_0/v_out_nand vdd fulladder_2/halfadder_0/nand_4/w_0_3# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1120 fulladder_2/halfadder_0/nand_0/a_13_n14# b3_4bitadder gnd Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1121 fulladder_2/halfadder_0/nand_0/v_out_nand a3_4bitadder fulladder_2/halfadder_0/nand_0/a_13_n14# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1122 fulladder_2/halfadder_0/nand_0/v_out_nand b3_4bitadder vdd fulladder_2/halfadder_0/nand_0/w_0_3# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1123 fulladder_2/halfadder_0/nand_0/v_out_nand a3_4bitadder vdd fulladder_2/halfadder_0/nand_0/w_0_3# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1124 fulladder_2/halfadder_0/nand_1/a_13_n14# fulladder_2/halfadder_0/nand_0/v_out_nand gnd Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1125 fulladder_2/halfadder_0/nand_1/v_out_nand b3_4bitadder fulladder_2/halfadder_0/nand_1/a_13_n14# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1126 fulladder_2/halfadder_0/nand_1/v_out_nand fulladder_2/halfadder_0/nand_0/v_out_nand vdd fulladder_2/halfadder_0/nand_1/w_0_3# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1127 fulladder_2/halfadder_0/nand_1/v_out_nand b3_4bitadder vdd fulladder_2/halfadder_0/nand_1/w_0_3# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1128 fulladder_2/halfadder_0/nand_2/a_13_n14# fulladder_2/halfadder_0/nand_0/v_out_nand gnd Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1129 fulladder_2/halfadder_0/nand_2/v_out_nand a3_4bitadder fulladder_2/halfadder_0/nand_2/a_13_n14# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1130 fulladder_2/halfadder_0/nand_2/v_out_nand fulladder_2/halfadder_0/nand_0/v_out_nand vdd fulladder_2/halfadder_0/nand_2/w_0_3# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1131 fulladder_2/halfadder_0/nand_2/v_out_nand a3_4bitadder vdd fulladder_2/halfadder_0/nand_2/w_0_3# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1132 fulladder_2/halfadder_1/nand_3/a_13_n14# fulladder_2/halfadder_1/nand_1/v_out_nand gnd Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1133 s3_4bitadder fulladder_2/halfadder_1/nand_2/v_out_nand fulladder_2/halfadder_1/nand_3/a_13_n14# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1134 s3_4bitadder fulladder_2/halfadder_1/nand_1/v_out_nand vdd fulladder_2/halfadder_1/nand_3/w_0_3# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1135 s3_4bitadder fulladder_2/halfadder_1/nand_2/v_out_nand vdd fulladder_2/halfadder_1/nand_3/w_0_3# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1136 fulladder_2/halfadder_1/nand_4/a_13_n14# fulladder_2/halfadder_1/nand_0/v_out_nand gnd Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1137 fulladder_2/or_0/v_a_or fulladder_2/halfadder_1/nand_0/v_out_nand fulladder_2/halfadder_1/nand_4/a_13_n14# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1138 fulladder_2/or_0/v_a_or fulladder_2/halfadder_1/nand_0/v_out_nand vdd fulladder_2/halfadder_1/nand_4/w_0_3# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1139 fulladder_2/or_0/v_a_or fulladder_2/halfadder_1/nand_0/v_out_nand vdd fulladder_2/halfadder_1/nand_4/w_0_3# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1140 fulladder_2/halfadder_1/nand_0/a_13_n14# fulladder_2/halfadder_1/v_a_halfadder gnd Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1141 fulladder_2/halfadder_1/nand_0/v_out_nand fulladder_2/c_in_fulladder fulladder_2/halfadder_1/nand_0/a_13_n14# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1142 fulladder_2/halfadder_1/nand_0/v_out_nand fulladder_2/halfadder_1/v_a_halfadder vdd fulladder_2/halfadder_1/nand_0/w_0_3# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1143 fulladder_2/halfadder_1/nand_0/v_out_nand fulladder_2/c_in_fulladder vdd fulladder_2/halfadder_1/nand_0/w_0_3# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1144 fulladder_2/halfadder_1/nand_1/a_13_n14# fulladder_2/halfadder_1/nand_0/v_out_nand gnd Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1145 fulladder_2/halfadder_1/nand_1/v_out_nand fulladder_2/halfadder_1/v_a_halfadder fulladder_2/halfadder_1/nand_1/a_13_n14# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1146 fulladder_2/halfadder_1/nand_1/v_out_nand fulladder_2/halfadder_1/nand_0/v_out_nand vdd fulladder_2/halfadder_1/nand_1/w_0_3# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1147 fulladder_2/halfadder_1/nand_1/v_out_nand fulladder_2/halfadder_1/v_a_halfadder vdd fulladder_2/halfadder_1/nand_1/w_0_3# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1148 fulladder_2/halfadder_1/nand_2/a_13_n14# fulladder_2/halfadder_1/nand_0/v_out_nand gnd Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1149 fulladder_2/halfadder_1/nand_2/v_out_nand fulladder_2/c_in_fulladder fulladder_2/halfadder_1/nand_2/a_13_n14# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1150 fulladder_2/halfadder_1/nand_2/v_out_nand fulladder_2/halfadder_1/nand_0/v_out_nand vdd fulladder_2/halfadder_1/nand_2/w_0_3# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1151 fulladder_2/halfadder_1/nand_2/v_out_nand fulladder_2/c_in_fulladder vdd fulladder_2/halfadder_1/nand_2/w_0_3# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1152 fulladder_2/or_0/a_n15_n30# fulladder_2/or_0/v_b_or gnd Gnd nfet w=12 l=3
+  ad=156 pd=74 as=0 ps=0
M1153 fulladder_2/or_0/a_n15_n30# fulladder_2/or_0/v_a_or gnd Gnd nfet w=12 l=3
+  ad=0 pd=0 as=0 ps=0
M1154 c_4bitadder fulladder_2/or_0/a_n15_n30# gnd Gnd nfet w=16 l=3
+  ad=84 pd=44 as=0 ps=0
M1155 fulladder_2/or_0/a_n15_10# fulladder_2/or_0/v_a_or vdd fulladder_2/or_0/w_n32_2# pfet w=12 l=3
+  ad=156 pd=74 as=0 ps=0
M1156 vdd fulladder_2/or_0/a_n15_n30# c_4bitadder fulladder_2/or_0/w_78_2# pfet w=16 l=3
+  ad=0 pd=0 as=80 ps=42
M1157 fulladder_2/or_0/a_n15_n30# fulladder_2/or_0/v_b_or fulladder_2/or_0/a_n15_10# fulladder_2/or_0/w_n32_2# pfet w=12 l=3
+  ad=72 pd=36 as=0 ps=0
C0 b3_4bitadder fulladder_2/halfadder_0/nand_1/w_0_3# 2.46fF
C1 halfadder_0/nand_3/w_0_3# halfadder_0/nand_1/v_out_nand 2.46fF
C2 fulladder_1/halfadder_1/nand_0/v_out_nand fulladder_1/halfadder_1/nand_1/w_0_3# 2.46fF
C3 a3_4bitadder fulladder_2/c_in_fulladder 5.40fF
C4 b3_4bitadder fulladder_2/c_in_fulladder 5.76fF
C5 fulladder_1/halfadder_1/nand_4/w_0_3# vdd 2.26fF
C6 fulladder_1/halfadder_1/nand_0/w_0_3# vdd 2.26fF
C7 fulladder_1/or_0/v_b_or s2_4bitadder 3.60fF
C8 halfadder_0/nand_4/w_0_3# halfadder_0/nand_0/v_out_nand 4.92fF
C9 fulladder_1/halfadder_1/nand_3/w_0_3# vdd 2.26fF
C10 s3_4bitadder fulladder_2/or_0/v_b_or 3.78fF
C11 fulladder_0/halfadder_0/nand_0/w_0_3# vdd 2.26fF
C12 fulladder_2/halfadder_0/nand_0/v_out_nand fulladder_2/halfadder_0/nand_2/w_0_3# 2.46fF
C13 fulladder_2/halfadder_1/nand_3/w_0_3# fulladder_2/halfadder_1/nand_2/v_out_nand 2.46fF
C14 fulladder_1/halfadder_1/nand_2/w_0_3# vdd 2.26fF
C15 fulladder_0/halfadder_0/nand_2/w_0_3# fulladder_0/halfadder_0/nand_0/v_out_nand 2.46fF
C16 fulladder_2/halfadder_0/nand_0/w_0_3# a3_4bitadder 6.51fF
C17 halfadder_0/nand_0/v_out_nand halfadder_0/nand_2/w_0_3# 2.46fF
C18 b3_4bitadder fulladder_2/halfadder_0/nand_0/w_0_3# 2.46fF
C19 b2_4bitadder fulladder_1/halfadder_0/nand_2/w_0_3# 2.46fF
C20 fulladder_2/or_0/v_b_or fulladder_2/or_0/w_n32_2# 5.19fF
C21 halfadder_0/nand_0/w_0_3# a0_4bitadder 6.51fF
C22 fulladder_1/halfadder_1/nand_1/w_0_3# fulladder_1/halfadder_1/v_a_halfadder 2.46fF
C23 s1_4bitadder fulladder_0/or_0/v_b_or 3.42fF
C24 halfadder_0/nand_3/w_0_3# halfadder_0/nand_2/v_out_nand 2.46fF
C25 fulladder_2/halfadder_0/nand_1/w_0_3# vdd 2.26fF
C26 fulladder_0/halfadder_0/nand_2/w_0_3# vdd 2.26fF
C27 fulladder_2/halfadder_1/nand_3/w_0_3# vdd 2.26fF
C28 gnd b1_4bitadder 3.54fF
C29 fulladder_0/halfadder_0/nand_1/v_out_nand fulladder_0/halfadder_0/nand_3/w_0_3# 2.46fF
C30 fulladder_2/c_in_fulladder vdd 2.60fF
C31 a3_4bitadder gnd 7.25fF
C32 vdd fulladder_0/halfadder_0/nand_3/w_0_3# 2.26fF
C33 fulladder_2/halfadder_1/nand_0/w_0_3# fulladder_2/c_in_fulladder 6.51fF
C34 b3_4bitadder gnd 7.72fF
C35 fulladder_0/halfadder_1/nand_0/w_0_3# fulladder_0/halfadder_1/v_a_halfadder 2.46fF
C36 fulladder_0/c_in_fulladder fulladder_0/halfadder_1/nand_2/w_0_3# 2.46fF
C37 fulladder_0/halfadder_1/v_a_halfadder fulladder_0/halfadder_1/nand_1/w_0_3# 2.46fF
C38 fulladder_0/or_0/w_78_2# fulladder_0/or_0/a_n15_n30# 5.74fF
C39 fulladder_0/or_0/v_a_or fulladder_0/or_0/w_n32_2# 5.19fF
C40 halfadder_0/nand_4/w_0_3# vdd 2.26fF
C41 fulladder_1/halfadder_0/nand_0/v_out_nand fulladder_1/halfadder_0/nand_2/w_0_3# 2.46fF
C42 fulladder_1/halfadder_1/nand_2/v_out_nand fulladder_1/halfadder_1/nand_3/w_0_3# 2.46fF
C43 fulladder_2/halfadder_1/nand_2/w_0_3# vdd 2.26fF
C44 fulladder_2/halfadder_0/nand_4/w_0_3# vdd 2.26fF
C45 b3_4bitadder a3_4bitadder 10.80fF
C46 fulladder_2/halfadder_0/nand_0/w_0_3# vdd 2.26fF
C47 fulladder_0/halfadder_1/nand_2/w_0_3# vdd 2.26fF
C48 fulladder_2/halfadder_1/nand_2/w_0_3# fulladder_2/halfadder_1/nand_0/v_out_nand 2.46fF
C49 fulladder_2/halfadder_1/nand_3/w_0_3# fulladder_2/halfadder_1/nand_1/v_out_nand 2.46fF
C50 halfadder_0/nand_2/w_0_3# vdd 2.26fF
C51 fulladder_0/halfadder_0/nand_1/w_0_3# b1_4bitadder 2.46fF
C52 halfadder_0/nand_3/w_0_3# vdd 2.26fF
C53 fulladder_0/c_in_fulladder b1_4bitadder 12.60fF
C54 fulladder_1/or_0/a_n15_n30# fulladder_1/or_0/w_78_2# 5.74fF
C55 fulladder_0/or_0/w_n32_2# fulladder_0/or_0/v_b_or 5.19fF
C56 fulladder_1/halfadder_1/nand_0/v_out_nand fulladder_1/halfadder_1/nand_4/w_0_3# 4.92fF
C57 fulladder_0/halfadder_0/nand_4/w_0_3# fulladder_0/halfadder_0/nand_0/v_out_nand 4.92fF
C58 gnd s2_4bitadder 5.67fF
C59 fulladder_0/halfadder_1/nand_0/v_out_nand fulladder_0/halfadder_1/nand_2/w_0_3# 2.46fF
C60 b1_4bitadder vdd 8.22fF
C61 vdd fulladder_1/halfadder_0/nand_4/w_0_3# 2.26fF
C62 gnd s0_4bitadder 2.70fF
C63 fulladder_0/c_in_fulladder fulladder_0/halfadder_1/nand_0/w_0_3# 6.51fF
C64 fulladder_0/or_0/w_n32_2# fulladder_0/or_0/a_n15_10# 3.38fF
C65 fulladder_0/halfadder_1/nand_3/w_0_3# vdd 2.26fF
C66 fulladder_0/halfadder_0/nand_4/w_0_3# vdd 2.26fF
C67 fulladder_1/halfadder_1/nand_0/v_out_nand fulladder_1/halfadder_1/nand_2/w_0_3# 2.46fF
C68 fulladder_0/halfadder_1/nand_1/v_out_nand fulladder_0/halfadder_1/nand_3/w_0_3# 2.46fF
C69 fulladder_2/halfadder_0/nand_1/w_0_3# fulladder_2/halfadder_0/nand_0/v_out_nand 2.46fF
C70 a3_4bitadder vdd 7.77fF
C71 vdd fulladder_1/halfadder_0/nand_1/w_0_3# 2.26fF
C72 b3_4bitadder vdd 7.20fF
C73 s3_4bitadder gnd 2.52fF
C74 a3_4bitadder fulladder_2/halfadder_0/nand_2/w_0_3# 2.46fF
C75 fulladder_0/halfadder_1/nand_0/w_0_3# vdd 2.26fF
C76 fulladder_0/halfadder_0/nand_1/w_0_3# fulladder_0/halfadder_0/nand_0/v_out_nand 2.46fF
C77 gnd s1_4bitadder 2.52fF
C78 fulladder_1/c_in_fulladder vdd 2.60fF
C79 halfadder_0/nand_1/w_0_3# halfadder_0/nand_0/v_out_nand 2.46fF
C80 vdd fulladder_0/halfadder_1/nand_1/w_0_3# 2.26fF
C81 fulladder_1/halfadder_0/nand_0/w_0_3# vdd 2.26fF
C82 fulladder_1/or_0/a_n15_10# fulladder_1/or_0/w_n32_2# 3.38fF
C83 fulladder_1/or_0/w_n32_2# fulladder_1/or_0/v_b_or 5.19fF
C84 fulladder_1/halfadder_1/nand_0/w_0_3# fulladder_1/halfadder_1/v_a_halfadder 2.46fF
C85 fulladder_0/halfadder_0/nand_1/w_0_3# vdd 2.26fF
C86 fulladder_0/c_in_fulladder vdd 2.60fF
C87 fulladder_1/halfadder_1/nand_1/w_0_3# vdd 2.26fF
C88 b2_4bitadder gnd 8.67fF
C89 fulladder_1/halfadder_0/nand_2/v_out_nand fulladder_1/halfadder_0/nand_3/w_0_3# 2.46fF
C90 fulladder_2/halfadder_0/nand_4/w_0_3# fulladder_2/halfadder_0/nand_0/v_out_nand 4.92fF
C91 fulladder_0/c_in_fulladder s0_4bitadder 2.70fF
C92 fulladder_2/halfadder_0/nand_1/v_out_nand fulladder_2/halfadder_0/nand_3/w_0_3# 2.46fF
C93 vdd fulladder_1/halfadder_0/nand_3/w_0_3# 2.26fF
C94 fulladder_0/halfadder_1/nand_0/v_out_nand fulladder_0/halfadder_1/nand_1/w_0_3# 2.46fF
C95 fulladder_2/or_0/v_a_or fulladder_2/or_0/w_n32_2# 5.19fF
C96 fulladder_0/halfadder_1/nand_4/w_0_3# vdd 2.26fF
C97 b2_4bitadder fulladder_1/halfadder_0/nand_1/w_0_3# 2.46fF
C98 halfadder_0/nand_2/w_0_3# a0_4bitadder 2.46fF
C99 fulladder_2/halfadder_1/nand_0/w_0_3# vdd 2.26fF
C100 vdd s2_4bitadder 3.46fF
C101 fulladder_2/halfadder_0/nand_3/w_0_3# vdd 2.26fF
C102 fulladder_0/halfadder_1/nand_2/v_out_nand fulladder_0/halfadder_1/nand_3/w_0_3# 2.46fF
C103 fulladder_1/or_0/w_n32_2# fulladder_1/or_0/v_a_or 5.19fF
C104 s0_4bitadder vdd 3.78fF
C105 fulladder_2/halfadder_0/nand_2/w_0_3# vdd 2.26fF
C106 fulladder_1/c_in_fulladder b2_4bitadder 8.64fF
C107 b2_4bitadder fulladder_1/halfadder_0/nand_0/w_0_3# 8.97fF
C108 fulladder_1/halfadder_0/nand_0/v_out_nand fulladder_1/halfadder_0/nand_4/w_0_3# 4.92fF
C109 fulladder_1/halfadder_1/nand_1/v_out_nand fulladder_1/halfadder_1/nand_3/w_0_3# 2.46fF
C110 halfadder_0/nand_1/w_0_3# vdd 2.26fF
C111 fulladder_2/halfadder_1/nand_4/w_0_3# vdd 2.26fF
C112 halfadder_0/nand_1/w_0_3# b0_4bitadder 2.46fF
C113 fulladder_2/halfadder_1/nand_1/w_0_3# vdd 2.26fF
C114 fulladder_0/halfadder_1/nand_0/v_out_nand fulladder_0/halfadder_1/nand_4/w_0_3# 4.92fF
C115 s3_4bitadder vdd 3.92fF
C116 fulladder_2/halfadder_1/nand_0/w_0_3# fulladder_2/halfadder_1/v_a_halfadder 2.46fF
C117 fulladder_1/halfadder_0/nand_0/v_out_nand fulladder_1/halfadder_0/nand_1/w_0_3# 2.46fF
C118 halfadder_0/nand_0/w_0_3# vdd 2.26fF
C119 fulladder_0/halfadder_0/nand_0/w_0_3# b1_4bitadder 8.97fF
C120 s1_4bitadder vdd 3.92fF
C121 fulladder_2/halfadder_1/nand_2/w_0_3# fulladder_2/c_in_fulladder 2.46fF
C122 fulladder_2/halfadder_1/nand_4/w_0_3# fulladder_2/halfadder_1/nand_0/v_out_nand 4.92fF
C123 halfadder_0/nand_0/w_0_3# b0_4bitadder 2.46fF
C124 fulladder_2/halfadder_1/nand_1/w_0_3# fulladder_2/halfadder_1/nand_0/v_out_nand 2.46fF
C125 b2_4bitadder vdd 11.82fF
C126 fulladder_2/halfadder_0/nand_3/w_0_3# fulladder_2/halfadder_0/nand_2/v_out_nand 2.46fF
C127 fulladder_2/halfadder_1/nand_1/w_0_3# fulladder_2/halfadder_1/v_a_halfadder 2.46fF
C128 fulladder_1/c_in_fulladder fulladder_1/halfadder_1/nand_0/w_0_3# 6.51fF
C129 fulladder_2/or_0/a_n15_n30# fulladder_2/or_0/w_78_2# 5.74fF
C130 fulladder_0/halfadder_0/nand_2/v_out_nand fulladder_0/halfadder_0/nand_3/w_0_3# 2.46fF
C131 fulladder_0/halfadder_0/nand_2/w_0_3# b1_4bitadder 2.46fF
C132 fulladder_1/halfadder_0/nand_2/w_0_3# vdd 2.26fF
C133 fulladder_1/c_in_fulladder fulladder_1/halfadder_1/nand_2/w_0_3# 2.46fF
C134 fulladder_1/halfadder_0/nand_1/v_out_nand fulladder_1/halfadder_0/nand_3/w_0_3# 2.46fF
C135 fulladder_2/or_0/a_n15_10# fulladder_2/or_0/w_n32_2# 3.38fF
C136 c_4bitadder Gnd 228.11fF
C137 fulladder_2/or_0/a_n15_n30# Gnd 59.49fF
C138 fulladder_2/halfadder_1/nand_0/v_out_nand Gnd 106.15fF
C139 fulladder_2/c_in_fulladder Gnd 92.45fF
C140 fulladder_2/halfadder_1/nand_2/a_13_n14# Gnd 2.44fF
C141 fulladder_2/halfadder_1/nand_2/v_out_nand Gnd 43.65fF
C142 fulladder_2/halfadder_1/nand_1/a_13_n14# Gnd 2.44fF
C143 fulladder_2/halfadder_1/nand_1/v_out_nand Gnd 27.54fF
C144 fulladder_2/halfadder_1/nand_0/a_13_n14# Gnd 2.44fF
C145 fulladder_2/halfadder_1/v_a_halfadder Gnd 113.23fF
C146 fulladder_2/halfadder_1/nand_4/a_13_n14# Gnd 2.44fF
C147 fulladder_2/or_0/v_a_or Gnd 39.01fF
C148 fulladder_2/halfadder_1/nand_3/a_13_n14# Gnd 2.44fF
C149 s3_4bitadder Gnd 273.68fF
C150 fulladder_2/halfadder_0/nand_0/v_out_nand Gnd 106.15fF
C151 a3_4bitadder Gnd 863.14fF
C152 fulladder_2/halfadder_0/nand_2/a_13_n14# Gnd 2.44fF
C153 fulladder_2/halfadder_0/nand_2/v_out_nand Gnd 43.65fF
C154 fulladder_2/halfadder_0/nand_1/a_13_n14# Gnd 2.44fF
C155 fulladder_2/halfadder_0/nand_1/v_out_nand Gnd 27.54fF
C156 fulladder_2/halfadder_0/nand_0/a_13_n14# Gnd 2.44fF
C157 b3_4bitadder Gnd 827.77fF
C158 fulladder_2/halfadder_0/nand_4/a_13_n14# Gnd 2.44fF
C159 fulladder_2/or_0/v_b_or Gnd 69.28fF
C160 fulladder_2/halfadder_0/nand_3/a_13_n14# Gnd 2.44fF
C161 fulladder_1/or_0/a_n15_n30# Gnd 59.49fF
C162 fulladder_1/halfadder_1/nand_0/v_out_nand Gnd 106.15fF
C163 fulladder_1/c_in_fulladder Gnd 88.31fF
C164 fulladder_1/halfadder_1/nand_2/a_13_n14# Gnd 2.44fF
C165 fulladder_1/halfadder_1/nand_2/v_out_nand Gnd 43.65fF
C166 fulladder_1/halfadder_1/nand_1/a_13_n14# Gnd 2.44fF
C167 fulladder_1/halfadder_1/nand_1/v_out_nand Gnd 27.54fF
C168 fulladder_1/halfadder_1/nand_0/a_13_n14# Gnd 2.44fF
C169 fulladder_1/halfadder_1/v_a_halfadder Gnd 113.23fF
C170 fulladder_1/halfadder_1/nand_4/a_13_n14# Gnd 2.44fF
C171 fulladder_1/or_0/v_a_or Gnd 39.01fF
C172 fulladder_1/halfadder_1/nand_3/a_13_n14# Gnd 2.44fF
C173 s2_4bitadder Gnd 308.54fF
C174 fulladder_1/halfadder_0/nand_0/v_out_nand Gnd 106.15fF
C175 b2_4bitadder Gnd 1266.42fF
C176 fulladder_1/halfadder_0/nand_2/a_13_n14# Gnd 2.44fF
C177 fulladder_1/halfadder_0/nand_2/v_out_nand Gnd 43.65fF
C178 fulladder_1/halfadder_0/nand_1/a_13_n14# Gnd 2.44fF
C179 fulladder_1/halfadder_0/nand_1/v_out_nand Gnd 27.54fF
C180 fulladder_1/halfadder_0/nand_0/a_13_n14# Gnd 2.44fF
C181 fulladder_1/halfadder_0/nand_4/a_13_n14# Gnd 2.44fF
C182 fulladder_1/or_0/v_b_or Gnd 69.28fF
C183 fulladder_1/halfadder_0/nand_3/a_13_n14# Gnd 2.44fF
C184 fulladder_0/or_0/a_n15_n30# Gnd 59.49fF
C185 fulladder_0/halfadder_1/nand_0/v_out_nand Gnd 106.15fF
C186 fulladder_0/c_in_fulladder Gnd 87.98fF
C187 fulladder_0/halfadder_1/nand_2/a_13_n14# Gnd 2.44fF
C188 fulladder_0/halfadder_1/nand_2/v_out_nand Gnd 43.65fF
C189 fulladder_0/halfadder_1/nand_1/a_13_n14# Gnd 2.44fF
C190 fulladder_0/halfadder_1/nand_1/v_out_nand Gnd 27.54fF
C191 fulladder_0/halfadder_1/nand_0/a_13_n14# Gnd 2.44fF
C192 fulladder_0/halfadder_1/v_a_halfadder Gnd 113.23fF
C193 fulladder_0/halfadder_1/nand_4/a_13_n14# Gnd 2.44fF
C194 fulladder_0/or_0/v_a_or Gnd 39.01fF
C195 fulladder_0/halfadder_1/nand_3/a_13_n14# Gnd 2.44fF
C196 s1_4bitadder Gnd 294.18fF
C197 fulladder_0/halfadder_0/nand_0/v_out_nand Gnd 106.15fF
C198 b1_4bitadder Gnd 938.49fF
C199 fulladder_0/halfadder_0/nand_2/a_13_n14# Gnd 2.44fF
C200 fulladder_0/halfadder_0/nand_2/v_out_nand Gnd 43.65fF
C201 fulladder_0/halfadder_0/nand_1/a_13_n14# Gnd 2.44fF
C202 gnd Gnd 2147.71fF
C203 fulladder_0/halfadder_0/nand_1/v_out_nand Gnd 27.54fF
C204 fulladder_0/halfadder_0/nand_0/a_13_n14# Gnd 2.44fF
C205 fulladder_0/halfadder_0/nand_4/a_13_n14# Gnd 2.44fF
C206 fulladder_0/or_0/v_b_or Gnd 69.28fF
C207 vdd Gnd 1409.30fF
C208 fulladder_0/halfadder_0/nand_3/a_13_n14# Gnd 2.44fF
C209 halfadder_0/nand_0/v_out_nand Gnd 106.15fF
C210 halfadder_0/nand_2/a_13_n14# Gnd 2.44fF
C211 halfadder_0/nand_2/v_out_nand Gnd 43.65fF
C212 halfadder_0/nand_1/a_13_n14# Gnd 2.44fF
C213 halfadder_0/nand_1/v_out_nand Gnd 27.54fF
C214 halfadder_0/nand_0/a_13_n14# Gnd 2.44fF
C215 b0_4bitadder Gnd 58.77fF
C216 halfadder_0/nand_4/a_13_n14# Gnd 2.44fF
C217 halfadder_0/nand_3/a_13_n14# Gnd 2.44fF
C218 s0_4bitadder Gnd 359.90fF
